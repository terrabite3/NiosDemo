// QsysDemo.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module QsysDemo (
		inout  wire [7:0]  character_lcd_cond_DATA, // character_lcd_cond.DATA
		output wire        character_lcd_cond_ON,   //                   .ON
		output wire        character_lcd_cond_BLON, //                   .BLON
		output wire        character_lcd_cond_EN,   //                   .EN
		output wire        character_lcd_cond_RS,   //                   .RS
		output wire        character_lcd_cond_RW,   //                   .RW
		input  wire        clk_clk,                 //                clk.clk
		input  wire [3:0]  key_cond_export,         //           key_cond.export
		output wire [8:0]  ledg_cond_export,        //          ledg_cond.export
		output wire [17:0] ledr_cond_export,        //          ledr_cond.export
		input  wire        reset_reset_n,           //              reset.reset_n
		output wire [31:0] seven_seg_cond_export,   //     seven_seg_cond.export
		input  wire [17:0] sw_cond_export           //            sw_cond.export
	);

	wire  [31:0] cpu_data_master_readdata;                                     // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                  // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                  // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [16:0] cpu_data_master_address;                                      // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                   // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                         // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                        // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                    // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                              // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                           // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [16:0] cpu_instruction_master_address;                               // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                  // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_character_lcd_avalon_lcd_slave_chipselect;  // mm_interconnect_0:character_lcd_avalon_lcd_slave_chipselect -> character_lcd:chipselect
	wire   [7:0] mm_interconnect_0_character_lcd_avalon_lcd_slave_readdata;    // character_lcd:readdata -> mm_interconnect_0:character_lcd_avalon_lcd_slave_readdata
	wire         mm_interconnect_0_character_lcd_avalon_lcd_slave_waitrequest; // character_lcd:waitrequest -> mm_interconnect_0:character_lcd_avalon_lcd_slave_waitrequest
	wire   [0:0] mm_interconnect_0_character_lcd_avalon_lcd_slave_address;     // mm_interconnect_0:character_lcd_avalon_lcd_slave_address -> character_lcd:address
	wire         mm_interconnect_0_character_lcd_avalon_lcd_slave_read;        // mm_interconnect_0:character_lcd_avalon_lcd_slave_read -> character_lcd:read
	wire         mm_interconnect_0_character_lcd_avalon_lcd_slave_write;       // mm_interconnect_0:character_lcd_avalon_lcd_slave_write -> character_lcd:write
	wire   [7:0] mm_interconnect_0_character_lcd_avalon_lcd_slave_writedata;   // mm_interconnect_0:character_lcd_avalon_lcd_slave_writedata -> character_lcd:writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;               // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;               // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;            // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;            // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                   // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;             // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                  // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;              // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_nios_ram_s1_chipselect;                     // mm_interconnect_0:nios_ram_s1_chipselect -> nios_ram:chipselect
	wire  [31:0] mm_interconnect_0_nios_ram_s1_readdata;                       // nios_ram:readdata -> mm_interconnect_0:nios_ram_s1_readdata
	wire  [12:0] mm_interconnect_0_nios_ram_s1_address;                        // mm_interconnect_0:nios_ram_s1_address -> nios_ram:address
	wire   [3:0] mm_interconnect_0_nios_ram_s1_byteenable;                     // mm_interconnect_0:nios_ram_s1_byteenable -> nios_ram:byteenable
	wire         mm_interconnect_0_nios_ram_s1_write;                          // mm_interconnect_0:nios_ram_s1_write -> nios_ram:write
	wire  [31:0] mm_interconnect_0_nios_ram_s1_writedata;                      // mm_interconnect_0:nios_ram_s1_writedata -> nios_ram:writedata
	wire         mm_interconnect_0_nios_ram_s1_clken;                          // mm_interconnect_0:nios_ram_s1_clken -> nios_ram:clken
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                  // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                   // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                     // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                 // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_seven_seg_s1_chipselect;                    // mm_interconnect_0:seven_seg_s1_chipselect -> seven_seg:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_s1_readdata;                      // seven_seg:readdata -> mm_interconnect_0:seven_seg_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_s1_address;                       // mm_interconnect_0:seven_seg_s1_address -> seven_seg:address
	wire         mm_interconnect_0_seven_seg_s1_write;                         // mm_interconnect_0:seven_seg_s1_write -> seven_seg:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_s1_writedata;                     // mm_interconnect_0:seven_seg_s1_writedata -> seven_seg:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                         // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                           // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                            // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                              // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                          // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                             // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                              // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_ledg_s1_chipselect;                         // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                           // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                            // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire         mm_interconnect_0_ledg_s1_write;                              // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                          // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                            // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                             // mm_interconnect_0:key_s1_address -> key:address
	wire         irq_mapper_receiver0_irq;                                     // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                                  // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [character_lcd:reset, cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, key:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, nios_ram:reset, rst_translator:in_reset, seven_seg:reset_n, sw:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [cpu:reset_req, nios_ram:reset_req, rst_translator:reset_req_in]

	QsysDemo_character_lcd character_lcd (
		.clk         (clk_clk),                                                      //                clk.clk
		.reset       (rst_controller_reset_out_reset),                               //              reset.reset
		.address     (mm_interconnect_0_character_lcd_avalon_lcd_slave_address),     //   avalon_lcd_slave.address
		.chipselect  (mm_interconnect_0_character_lcd_avalon_lcd_slave_chipselect),  //                   .chipselect
		.read        (mm_interconnect_0_character_lcd_avalon_lcd_slave_read),        //                   .read
		.write       (mm_interconnect_0_character_lcd_avalon_lcd_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_character_lcd_avalon_lcd_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_character_lcd_avalon_lcd_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_character_lcd_avalon_lcd_slave_waitrequest), //                   .waitrequest
		.LCD_DATA    (character_lcd_cond_DATA),                                      // external_interface.export
		.LCD_ON      (character_lcd_cond_ON),                                        //                   .export
		.LCD_BLON    (character_lcd_cond_BLON),                                      //                   .export
		.LCD_EN      (character_lcd_cond_EN),                                        //                   .export
		.LCD_RS      (character_lcd_cond_RS),                                        //                   .export
		.LCD_RW      (character_lcd_cond_RW)                                         //                   .export
	);

	QsysDemo_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	QsysDemo_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	QsysDemo_key key (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata), //                    .readdata
		.in_port  (key_cond_export)                    // external_connection.export
	);

	QsysDemo_ledg ledg (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_cond_export)                      // external_connection.export
	);

	QsysDemo_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_cond_export)                      // external_connection.export
	);

	QsysDemo_nios_ram nios_ram (
		.clk        (clk_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_nios_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_nios_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_nios_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_nios_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_nios_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_nios_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_nios_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)        //       .reset_req
	);

	QsysDemo_seven_seg seven_seg (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_cond_export)                      // external_connection.export
	);

	QsysDemo_sw sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_cond_export)                    // external_connection.export
	);

	QsysDemo_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                       //   irq.irq
	);

	QsysDemo_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	QsysDemo_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                (clk_clk),                                                      //                         clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                               // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                    (cpu_data_master_address),                                      //                 cpu_data_master.address
		.cpu_data_master_waitrequest                (cpu_data_master_waitrequest),                                  //                                .waitrequest
		.cpu_data_master_byteenable                 (cpu_data_master_byteenable),                                   //                                .byteenable
		.cpu_data_master_read                       (cpu_data_master_read),                                         //                                .read
		.cpu_data_master_readdata                   (cpu_data_master_readdata),                                     //                                .readdata
		.cpu_data_master_write                      (cpu_data_master_write),                                        //                                .write
		.cpu_data_master_writedata                  (cpu_data_master_writedata),                                    //                                .writedata
		.cpu_data_master_debugaccess                (cpu_data_master_debugaccess),                                  //                                .debugaccess
		.cpu_instruction_master_address             (cpu_instruction_master_address),                               //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest         (cpu_instruction_master_waitrequest),                           //                                .waitrequest
		.cpu_instruction_master_read                (cpu_instruction_master_read),                                  //                                .read
		.cpu_instruction_master_readdata            (cpu_instruction_master_readdata),                              //                                .readdata
		.character_lcd_avalon_lcd_slave_address     (mm_interconnect_0_character_lcd_avalon_lcd_slave_address),     //  character_lcd_avalon_lcd_slave.address
		.character_lcd_avalon_lcd_slave_write       (mm_interconnect_0_character_lcd_avalon_lcd_slave_write),       //                                .write
		.character_lcd_avalon_lcd_slave_read        (mm_interconnect_0_character_lcd_avalon_lcd_slave_read),        //                                .read
		.character_lcd_avalon_lcd_slave_readdata    (mm_interconnect_0_character_lcd_avalon_lcd_slave_readdata),    //                                .readdata
		.character_lcd_avalon_lcd_slave_writedata   (mm_interconnect_0_character_lcd_avalon_lcd_slave_writedata),   //                                .writedata
		.character_lcd_avalon_lcd_slave_waitrequest (mm_interconnect_0_character_lcd_avalon_lcd_slave_waitrequest), //                                .waitrequest
		.character_lcd_avalon_lcd_slave_chipselect  (mm_interconnect_0_character_lcd_avalon_lcd_slave_chipselect),  //                                .chipselect
		.cpu_debug_mem_slave_address                (mm_interconnect_0_cpu_debug_mem_slave_address),                //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                  (mm_interconnect_0_cpu_debug_mem_slave_write),                  //                                .write
		.cpu_debug_mem_slave_read                   (mm_interconnect_0_cpu_debug_mem_slave_read),                   //                                .read
		.cpu_debug_mem_slave_readdata               (mm_interconnect_0_cpu_debug_mem_slave_readdata),               //                                .readdata
		.cpu_debug_mem_slave_writedata              (mm_interconnect_0_cpu_debug_mem_slave_writedata),              //                                .writedata
		.cpu_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_debug_mem_slave_byteenable),             //                                .byteenable
		.cpu_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),            //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),            //                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                .write
		.jtag_uart_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                .read
		.jtag_uart_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                .chipselect
		.key_s1_address                             (mm_interconnect_0_key_s1_address),                             //                          key_s1.address
		.key_s1_readdata                            (mm_interconnect_0_key_s1_readdata),                            //                                .readdata
		.ledg_s1_address                            (mm_interconnect_0_ledg_s1_address),                            //                         ledg_s1.address
		.ledg_s1_write                              (mm_interconnect_0_ledg_s1_write),                              //                                .write
		.ledg_s1_readdata                           (mm_interconnect_0_ledg_s1_readdata),                           //                                .readdata
		.ledg_s1_writedata                          (mm_interconnect_0_ledg_s1_writedata),                          //                                .writedata
		.ledg_s1_chipselect                         (mm_interconnect_0_ledg_s1_chipselect),                         //                                .chipselect
		.ledr_s1_address                            (mm_interconnect_0_ledr_s1_address),                            //                         ledr_s1.address
		.ledr_s1_write                              (mm_interconnect_0_ledr_s1_write),                              //                                .write
		.ledr_s1_readdata                           (mm_interconnect_0_ledr_s1_readdata),                           //                                .readdata
		.ledr_s1_writedata                          (mm_interconnect_0_ledr_s1_writedata),                          //                                .writedata
		.ledr_s1_chipselect                         (mm_interconnect_0_ledr_s1_chipselect),                         //                                .chipselect
		.nios_ram_s1_address                        (mm_interconnect_0_nios_ram_s1_address),                        //                     nios_ram_s1.address
		.nios_ram_s1_write                          (mm_interconnect_0_nios_ram_s1_write),                          //                                .write
		.nios_ram_s1_readdata                       (mm_interconnect_0_nios_ram_s1_readdata),                       //                                .readdata
		.nios_ram_s1_writedata                      (mm_interconnect_0_nios_ram_s1_writedata),                      //                                .writedata
		.nios_ram_s1_byteenable                     (mm_interconnect_0_nios_ram_s1_byteenable),                     //                                .byteenable
		.nios_ram_s1_chipselect                     (mm_interconnect_0_nios_ram_s1_chipselect),                     //                                .chipselect
		.nios_ram_s1_clken                          (mm_interconnect_0_nios_ram_s1_clken),                          //                                .clken
		.seven_seg_s1_address                       (mm_interconnect_0_seven_seg_s1_address),                       //                    seven_seg_s1.address
		.seven_seg_s1_write                         (mm_interconnect_0_seven_seg_s1_write),                         //                                .write
		.seven_seg_s1_readdata                      (mm_interconnect_0_seven_seg_s1_readdata),                      //                                .readdata
		.seven_seg_s1_writedata                     (mm_interconnect_0_seven_seg_s1_writedata),                     //                                .writedata
		.seven_seg_s1_chipselect                    (mm_interconnect_0_seven_seg_s1_chipselect),                    //                                .chipselect
		.sw_s1_address                              (mm_interconnect_0_sw_s1_address),                              //                           sw_s1.address
		.sw_s1_readdata                             (mm_interconnect_0_sw_s1_readdata),                             //                                .readdata
		.sys_clk_timer_s1_address                   (mm_interconnect_0_sys_clk_timer_s1_address),                   //                sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                     (mm_interconnect_0_sys_clk_timer_s1_write),                     //                                .write
		.sys_clk_timer_s1_readdata                  (mm_interconnect_0_sys_clk_timer_s1_readdata),                  //                                .readdata
		.sys_clk_timer_s1_writedata                 (mm_interconnect_0_sys_clk_timer_s1_writedata),                 //                                .writedata
		.sys_clk_timer_s1_chipselect                (mm_interconnect_0_sys_clk_timer_s1_chipselect),                //                                .chipselect
		.sysid_control_slave_address                (mm_interconnect_0_sysid_control_slave_address),                //             sysid_control_slave.address
		.sysid_control_slave_readdata               (mm_interconnect_0_sysid_control_slave_readdata)                //                                .readdata
	);

	QsysDemo_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
